library verilog;
use verilog.vl_types.all;
entity REGISTRADOR_32BIT_vlg_vec_tst is
end REGISTRADOR_32BIT_vlg_vec_tst;
